  typedef struct{
  	integer rmode;
    integer fpu_op;
    shortreal opa;
    shortreal opb;
    shortreal resultado;
  } packet;